`timescale 1ns / 1ps

module InstructionMemory(
    input clk,
    input rsta,
    input [31:0]  addra,
    output [31:0] douta
);
    integer i;

	reg	[31:0]	IMem[0:127];	// A size of 128 instrutions each with size 32 bits.
	always @(posedge clk) begin
        if(rsta) begin
            	IMem[0] = 32'b00000110001101010000000000000000;
                IMem[1] = 32'b01000110001000000000000000000000;
                IMem[2] = 32'b00000110000000010000000000000001;
                IMem[3] = 32'b00100110001000100000000000000000;
                IMem[4] = 32'b00010100101001010000000000000000;
                IMem[5] = 32'b00010100001100000000000000000000;
                IMem[6] = 32'b00010110101101010000000000000000;
                IMem[7] = 32'b00010100000000000000000000000000;
                IMem[8] = 32'b01010100110000000000000000000001;
                IMem[9] = 32'b01010100110100000000000000000000;
                IMem[10] = 32'b00011100111001010000000000000000;
                IMem[11] = 32'b00011100110000000000000000000000;
                IMem[12] = 32'b00011110110100100000000000000000;
                IMem[13] = 32'b00011100111100000000000000000000;
                IMem[14] = 32'b11000000000001110000000000000100;
                IMem[15] = 32'b10010100110000000000000000000000;
                IMem[16] = 32'b10010100110100000000000000000001;
                IMem[17] = 32'b00010110101101010000000000000000;
                IMem[18] = 32'b00010110000000010000000000000001;
                IMem[19] = 32'b00010100000000010000000000000001;
                IMem[20] = 32'b00100001000001010000000000000000;
                IMem[21] = 32'b00100000101000000000000000000000;
                IMem[22] = 32'b00100001001100000000000000000000;
                IMem[23] = 32'b11000000000001101111111111101111;
                IMem[24] = 32'b00010110000000000000000000000000;
                IMem[25] = 32'b11000000000000111111111111101010;
                IMem[26] = 32'b01000111100100000000000000000000;
                IMem[27] = 32'b00110010000000000000000000000000;
                IMem[28] = 32'b00000110000000010000000000000001;
                IMem[29] = 32'b00000100000000011111111111111111;
                IMem[30] = 32'b11000000000000111111111111111011;
                IMem[31] = 32'b11000000000000111111111111111011;	
                for (i = 32; i < 128; i = i + 1) begin
                    IMem[i] = 32'b0;
                end 
        end  
	end
	 

	assign  douta = IMem[addra];


endmodule
